* Josephson junction component test
* Date modified: 2020/01/22
B1  1   0  jj1   area=1
Itest   0   1   pwl(0 0 10p 0 50p 250u 200p 250u 240p 0 250p 0 300p -250u 450p -250u 500p 0)
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.tran 0.01p 500p
.print devv B1
.print devi B1
.print devp B1