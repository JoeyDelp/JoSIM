* jj_pump.js
ISin    0          1          SIN(0 0.2mA 80GHz 200ps 0)
IDC 	0	   1	      PWL(0 0 10p 0 50p 2.5E-7)
B1      1          2          jj1        area=1
R1      1          2          8
RS	2	   0	      2        
.model jj1 jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rN=16, icrit=0.1mA)
.tran 0.05p 500p 0 0.25p
.print DEVI ISin
.print NODEV 1 0
.end
