Vin	1	0	pwl(0 0 50p 0 52p 5 55p 5 57p 0)
RL	1	2	20
T1	2	0	3	0	lossless TD=100p Z0=100
T2	3	0	4	0	lossless TD=100p Z0=100
T3	4	0	5	0	lossless TD=100p Z0=100
T4	5	0	6	0	lossless TD=100p Z0=100
T5	6	0	7	0	lossless TD=100p Z0=100
T6	7	0	8	0	lossless TD=100p Z0=100
T7	8	0	9	0	lossless TD=100p Z0=100
T8	9	0	10	0	lossless TD=100p Z0=100
Rout	10	0	20
.tran 0.25p 3000p 0 0.25p
.print nodev 1
.print nodev 2
.print nodev 3
.print nodev 4
.print nodev 5
.print nodev 6
.print nodev 7
.print nodev 8
.print nodev 9
.print nodev 10
.end
